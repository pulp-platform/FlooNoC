// Copyright 2024 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Lukas Berner <bernerl@student.ethz.ch>

// sa local: choose a valid vc via rr arbitration
module floo_look_ahead_routing #( )(
    input logic                 vc_ctrl_head_vld_i,
    input hdr_t                 vc_ctrl_head_i,

    output route_dir_e          look_ahead_routing_o,

    input id_t                  xy_id_i
);





endmodule
