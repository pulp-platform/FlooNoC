/*test ideas:
1) connectivity from each input vs to each output vc, lookahead is set correctly on output
2) FVADA working correctly: forward to different vc if prioritized one is not free -> lookahead still set correctly
3) dont send if all buffers full





*/