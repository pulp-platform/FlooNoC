// Copyright 2022 ETH Zurich and University of Bologna.
// Solderpad Hardware License, Version 0.51, see LICENSE for details.
// SPDX-License-Identifier: SHL-0.51
//
// Tim Fischer <fischeti@iis.ee.ethz.ch>

package floo_test_pkg;

  typedef enum {
    FastSlave,
    SlowSlave,
    MixedSlave
  } slave_type_e;

endpackage
